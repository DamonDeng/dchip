module tb;

initial begin
    $display("*************************");
    $display("hello world");
    $display("*************************");
end

endmodule

